// FP-UVM - UVM for FPGAs app 
// Automatically generated from VHDL Package: NUMERIC_STD 
package sv_NUMERIC_STD; 
  parameter CopyRightNotice = 256618540;
  parameter NAU = 256618540;
  parameter NAS = 256618540;
  parameter NO_WARNING = 0;
  parameter MATCH_TABLE = 0;
endpackage : sv_NUMERIC_STD 

import sv_NUMERIC_STD::* 

