// FP-UVM - UVM for FPGAs app 
// Automatically generated from VHDL Package: types_common 
package sv_types_common; 
  parameter log2 = 0;
  parameter log2x = 0;
  parameter zero32 = 0;
  parameter zero64 = 0;
endpackage : sv_types_common 

import sv_types_common::* 

