// FP-UVM - UVM for FPGAs app 
// Automatically generated from VHDL Package: gencomp 
package sv_gencomp; 
  parameter NTECH = 53;
  parameter inferred = 0;
  parameter virtex = 1;
  parameter virtex2 = 2;
  parameter memvirage = 3;
  parameter axcel = 4;
  parameter proasic = 5;
  parameter atc18s = 6;
  parameter altera = 7;
  parameter umc = 8;
  parameter rhumc = 9;
  parameter apa3 = 10;
  parameter spartan3 = 11;
  parameter ihp25 = 12;
  parameter rhlib18t = 13;
  parameter virtex4 = 14;
  parameter lattice = 15;
  parameter ut25 = 16;
  parameter spartan3e = 17;
  parameter peregrine = 18;
  parameter memartisan = 19;
  parameter virtex5 = 20;
  parameter custom1 = 21;
  parameter ihp25rh = 22;
  parameter stratix1 = 23;
  parameter stratix2 = 24;
  parameter eclipse = 25;
  parameter stratix3 = 26;
  parameter cyclone3 = 27;
  parameter memvirage90 = 28;
  parameter tsmc90 = 29;
  parameter easic90 = 30;
  parameter atc18rha = 31;
  parameter smic013 = 32;
  parameter tm65gpl = 33;
  parameter axdsp = 34;
  parameter spartan6 = 35;
  parameter virtex6 = 36;
  parameter actfus = 37;
  parameter stratix4 = 38;
  parameter st65lp = 39;
  parameter st65gp = 40;
  parameter easic45 = 41;
  parameter cmos9sf = 42;
  parameter apa3e = 43;
  parameter apa3l = 44;
  parameter ut130 = 45;
  parameter ut90 = 46;
  parameter gf65 = 47;
  parameter virtex7 = 48;
  parameter kintex7 = 49;
  parameter artix7 = 50;
  parameter zynq7000 = 51;
  parameter rhlib13t = 52;
  parameter mikron180 = 53;
  parameter is_fpga = 53;
endpackage : sv_gencomp 

import sv_gencomp::* 

