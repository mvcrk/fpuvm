// FP-UVM - UVM for FPGAs app 
// Automatically generated from VHDL Package: NUMERIC_STD 
package sv_NUMERIC_STD; 
  parameter CopyRightNotice = 1715212332;
  parameter NAU = 1715212332;
  parameter NAS = 1715212332;
  parameter NO_WARNING = 0;
  parameter MATCH_TABLE = 0;
endpackage : sv_NUMERIC_STD 

import sv_NUMERIC_STD::* 

